module Mux1(input logic In1, In2, Control, output logic Out);
	always_comb begin
		if(Control == 0)
			Out <= In1;
		else 
			Out <= In2;
	end

endmodule // mux